module elelock(key, lock);
    input key;
    output lock;
endmodule